grammar edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:sqliteOn;

exports edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:sqliteOn:query;

