grammar edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:foreach;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOnQuery;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOnCommit;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:types;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:use;


