grammar determinism;

import edu:umn:cs:melt:ableC:host;


copper_mda foreachStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:foreach;
}


copper_mda useStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:use;
}


copper_mda foreachStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:foreach;
}


copper_mda sqliteOnQuery(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:sqliteOnQuery;
}


copper_mda sqliteOnCommit(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:sqliteOnCommit;
}



