grammar edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax:foreach;
exports edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax:sqliteOn;
exports edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax:tables;
exports edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax:types;
exports edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax:use;

global builtin::Location = loc("Built In", 0, 0, 0, 0, 0, 0);
