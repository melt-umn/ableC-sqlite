grammar determinism;

import edu:umn:cs:melt:ableC:host;


copper_mda foreachStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:foreach;
}


copper_mda useStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:use;
}


copper_mda foreachStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:foreach;
}


copper_mda sqliteOnQuery(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOnQuery;
}


copper_mda sqliteOnCommit(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOnCommit;
}



