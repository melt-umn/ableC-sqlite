grammar edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:onKeyword;

imports edu:umn:cs:melt:ableC:concretesyntax;

marking terminal SqliteOn_t 'on' lexer classes {Ckeyword};
