grammar edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax:sqliteOn;

exports edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax:sqliteOn:query;
