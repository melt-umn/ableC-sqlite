grammar edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax:sqliteOn;

exports edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax:sqliteOn:query;
