grammar edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOn;

exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOn:query;

