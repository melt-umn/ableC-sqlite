grammar edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:foreach;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOn;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:types;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:use;

