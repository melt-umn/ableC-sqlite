grammar edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax:foreach;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax:sqliteOn;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax:tables;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax:types;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax:use;

