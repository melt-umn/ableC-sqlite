grammar edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:foreach;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:sqliteOnQuery;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:sqliteOnCommit;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:types;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax:use;


