grammar edu:umn:cs:melt:exts:ableC:sqlite:modular_analyses:determinism;

import edu:umn:cs:melt:ableC:host;

copper_mda testStmt(ablecParser) {
  edu:umn:cs:melt:ableC:host;
  edu:umn:cs:melt:exts:ableC:sqlite;
}

