grammar edu:umn:cs:melt:exts:ableC:sqlite:src;

exports edu:umn:cs:melt:exts:ableC:sqlite:src:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:sqlite:src:concretesyntax;

